----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 26.02.2021 09:22:36
-- Design Name: 
-- Module Name: Dec_3v8 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Dec_3v8 is
    Port ( E : in STD_LOGIC_VECTOR (2 downto 0);
           S : out STD_LOGIC_VECTOR (7 downto 0));
end Dec_3v8;

architecture Behavioral of Dec_3v8 is

begin

with E select
S <=    x"01" when "000",
        x"02" when "001",
        x"04" when "010",
        x"08" when "011",
        x"10" when "100",
        x"20" when "101",
        x"40" when "110",
        x"80" when "111",
        "--------" when others;
        
        
        

end Behavioral;
